13375||Aldenham|the county of Shropshire
13368|||
13369||Thornes|the county of West Yorkshire
13370||Rotherham|the county of South Yorkshire
13371||Knock|the city of Belfast
13381|Abbeydale|the city of Sheffield|
13105|Megiddo||
13104||Norbury|the London Borough of Croydon
13103|Liverpool|Mossley Hill|the county of Merseyside
13102||Brondesbury|the London Borough of Brent
13109|||
13108||Southover|the county of East Sussex
13107|St Johns||the county of Surrey
13106|Sandwell||the county of West Midlands
13097|Weston-super-Mare||
13096|Ilminster|Ashill|the county of Somerset
12883|Arran||
12884||Chichester|the county of West Sussex
10015|Norton-sub-Hamdon||the county of Somerset
12882|Stoke|Widnes|the county of Cheshire
12879|Upholland|St Albans|the county of Hertfordshire
12880|||
12877|Hever||
12878||Richmond upon Thames|the London Borough of Richmond upon Thames
12875|||
12876|||
13526||Lutterworth|the county of Leicestershire
13525||Regent's Park|the city of Westminster
13528|Dorking|Iford|the county of East Sussex
13527|Bewdley||
13521|Tewkesbury|Gotherington|the county of Gloucestershire
13524||Anagach|Highland
13523||Heywood and Royton|Greater Manchester
13512|Brighton||the county of East Sussex
13511|Whitley|Child's Hill|Greater London
13503||Belgravia|the city of Westminster
13505||Cranford|the London Borough of Hilllingdon
13506|Craigweil||the county of West Sussex
13507||Godmanstone|the county of Dorset
13508||Hampton|the London Borough of Richmond
13509||Tanat|the county of Shropshire
13510||Banbury|the county of Oxfordshire
13501|Cornhill|Boughrood|the county of Powys
13502||Liverpool|the county of Merseyside
13711|Crossharbour||the London Borough of Tower Hamlets
13241||Stoke Newington|Greater London
13240||Woodcote|the county of Surrey
13238||Blackpool|the county of Lancashire and of Lindfield in the County of West Sussex
13236||Cromac|the city of Belfast
13367|||
13692||Blackwatertown|the county of Armagh
12981|Rowington||the county of Warwickshire
10054||Sandwell|the county of West Midlands
12980||Abbots Morton|the county of Hereford and Worcester
12985|Faversham||the county of Kent
12986||Warlingham|the county of Surrey and of Croydon in the London Borough of Croydon
12983||Pimlico|the city of Westminster
12984|Tara||
13028||Wallingford|the county of Oxfordshire
13034||Wigton|the county of Cumbria
13636||Bushfield|the county of Hampshire
13635||Bibury|the county of Gloucestershire
13638||Lydd|the county of Kent
13637|Harwich||the county of Essex
13640|||
13639|||
13642||Lewes|the county of East Sussex
13610|Spennithorne||the county of North Yorkshire
13611|Alverthorpe||the county of West Yorkshire
10067|Sutton Mandeville||the county of Wiltshire
13613|||
13606||Ebbw Vale|the county of Gwent
13607|Tremorfa||the county of South Glamorgan
13608|||
13609|Madingley|Cambridge|the county of Cambridgeshire
13604||Camden|the London Borough of Camden
13343||Rowlands Gill|the county of Tyne and Wear
13430||Pitshanger|the London Borough of Ealing
13451||Goring|the county of Oxfordshire
13347|Brockwell|Herne Hill|the London Borough of Lambeth
13345|Alsa|Stiffkey|the county of Norfolk
13458||Rothley|the county of Leicestershire
13351|Caithness||
13676|Lochbroom||the District of Ross and Cromarty
13679|Alloway|Ayr|the District of Kyle and Carrick
10090||Allerdale|the county of Cumbria
13672|Canterbury||
13669|Clifton||the city and county of Bristol
13674|Berriew||the county of Powys
13670|Lour||the District of Angus
13018|Hadley|Monken Hadley|Greater London
13019||Upton|the county of Nottinghamshire
13016||Devizes|the county of Wiltshire
13017|Furness|Cartmel|the county of Cumbria
13014||Dean|the county of Oxfordshire
13015||Llantarnam|the county of Monmouth
13012|Wallasey|Leigh-on-Sea|the county of Essex
13010||Aldershot|the county of Hampshire
13253|Chester||
13252||Cranfield|the county of Bedfordshire
13251||Ryedale|the county of North Yorkshire
13258|Cholmondeley||
13257|||
13256||Leckhampton|the county of Gloucestershire
10108|Windermere||the county of Cumbria
13248|Hampstead||the London Borough of Camden
13517||Clapham|the London Borough of Lambeth
13518||Hackney|the London Borough of Hackney
13519||Briglands|Perthshire and Kinross
13520|||
13513||Dover|the county of Kent
13514||Ranmore|the county of Surrey
13515|Pimlico||the city of Westminster
13516|Culross||
13550|||
13556||Langton Green|the county of Kent
12869|Islandreagh||the county of Antrim
12872|Thorndon|Wellington|New Zealand and of Cambridge in the county of Cambridgeshire
12871|Berkeley||the county of Gloucestershire
10132|Castle Vale|Erdington|the county of West Midlands
12873|Courtown||
13585|Coventry||
13559||Queensbury|Greater London
13235|Radley|Helhoughton|the county of Norfolk
13599|||
12952|||
12954|Crawford and Balcarres||
13094||Edgbaston|the county of West Midlands
13095||Pont Esgob|the Black Mountains and the county of Powys
13100||the London Borough of Croydon|
13101||Millbank|the city of Westminster
13098|Whitekirk||East Lothian
13099||Newick|the county of East Sussex
12966|Marylebone||the city of Westminster
13399||Clare Market|the city of Westminster
13398|||
13397||Romsey|the city of Cambridge
13396|Coity|Penybont|the county of Mid Glamorgan
13395|Oldham|Broxbourne|the county of Hertfordshire
13394|Harptree|Wedmore|the county of Somerset
13393|Thornton-le-Fylde|Eccles|the county of Greater Manchester
13392||Kingston upon Hull|the county of the East Riding of Yorkshire
13391||Aldington|the county of Kent
13390|Alteryn||the county of Gwent
13659|||
13661||St Clement Danes|the city of Westminster
13662||Waltham Brooks|the county of West Sussex
13664||Jarrow|the county of Tyne and Wear
13665||Bocking|the county of Essex
13651||Ashton|the county of Northamptonshire
13000||Battersea|the London Borough of Wandsworth
12999|Dundee||
13002||Hong Kong Island|Hong Kong and of Knightsbridge in the Royal Borough of Kensington and Chelsea
12996|Durham||
12995||Armagh|the county of Armagh
12998||Stratton St Margaret|the county of Wiltshire
12997|Moulton||the county of North Yorkshire
13004|Winton|Rushyford|the county of Durham
13003||Kirkcaldy|Fife
13234||Nant Conwy|the county of Gwynedd
13696||the city of Westminster|
13232|Morpeth||the county of Northumberland and of the city of Newcastle upon Tyne
13233|||
13230||Aberteifi|the county of Dyfed
13231||Tunbridge Wells|the county of Kent and of Clerkenwell in the London Borough of Islington
13229|Erroll||
13242|Parkside|St Helens|the county of Merseyside
13243|Temple Guiting||the county of Gloucestershire
12852|Watford|Chipperfield|the county of Hertfordshire
12853|Kirkford|Cowdenbeath|the District of Dunfermline
12850||Horsham|the county of West Sussex
12851|Thoroton||the county of Nottinghamshire
12848||West Haddon|Northamptonshire
12849|Falkland||
12846|Ribbleton|Fulwood|the county of Lancashire
12847|Worcester|Wimbledon|the London Borough of Merton
10196||Southport|the county of Merseyside
12855||Frognal|the London Borough of Camden
13470||Shotesham|the county of Norfolk
13469|||
13472||Pimlico|the city of Westminster
13471|Llandaff||the county of South Glamorgan
13468|||
13467||Queen's Gate|the city of Westminster
13474||Plymouth|the county of Devon
13473|Drumlean||Stirling
13311||Ripley|the county of Surrey
13312|Thames Bank|Reddish|the county of Greater Manchester
10212||Sutton Coldfield|the county of West Midlands
13314|Carmyllie||the District of Angus
13307||Dingley|the county of Northamptonshire
13308|||
13309|Fairfield|Sauchie|the county of Clackmannanshire
13310||Blaenrhondda|the county of Mid Glamorgan
13304|Parkes|Southgate|Greater London and of Parkes in the State of New South Wales and Commonwealth of Australia
13063||Watford|the county of Hertfordshire
13062||Highgate|the London Borough of Camden
13061|||
13066|Market Rasen||the county of Lincolnshire
13065||Dudley|the county of West Midlands
13064|Craigmillar||the District of the city of Edinburgh
13068||Glenridding|the county of Cumbria
12919|||
12920|||
12918|Chieveley||the Royal county of Berkshire
10233||Newcastle-under-Lyme|the county of Staffordshire
12924||Allerton|the county of Merseyside
12921||Youlbury|the county of Oxfordshire
12922|Strathblane|Deil's Craig|Stirling
12914|||
12915||Roundwood|the London Borough of Brent
13569|Potternewton|Leeds|the county of West Yorkshire
13568||Aldwych|the city of Westminster
13571|Edmonton||Greater London
13570|||
13572||Pendle|the county of Lancashire
13574||Ot Moor|the county of Oxfordshire
13561||Notting Hill|the Royal Borough of Kensington and Chelsea
13560|||
13414||Stockport|Greater Manchester
13415||Kilvey|the county of Swansea
13416||Govilon|the county of Gwent
13417|Fforestfach||the county of West Glamorgan
10247||Telford|the county of Shropshire
13420|Craigiebank||the city of Dundee
13421||Calverton|the county of Buckinghamshire
13422||Richmond upon Thames|the London Borough of Richmond upon Thames
13423||Kensington|the Royal Borough of Kensington and Chelsea
13140|Chiswick|Bedford Park|the London Borough of Ealing
13139||Chelmsford|the county of Essex
13137||Blackford|the city of Edinburgh
13135|Haringey|Hornsey|the London Borough of Haringey
13134|High Cross|Tottenham|Greater London
13133|Peckham||the London Borough of Southwark
13148|Richmond||the county of North Yorkshire
13147||Chester|the county of Cheshire
13499||Higher Broughton|the county of Greater Manchester
13500||Skidby|the county of the East Riding of Yorkshire
13497||Sparkbrook|the county of West Midlands
13498||Isleworth|the London Borough of Hounslow
13495||Dartmouth Park|the London Borough of Camden
13496||Riddlesden|the county of West Yorkshire
13493|||
10276||Thenford|the county of Northamptonshire
13340||Worthing|the county of West Sussex
13224|Eggardon||the county of Dorset
13226|Astley Abbotts|Nash|the county of Shropshire
13221||Chedworth|the county of Gloucestershire
13220||Kettlethorpe|the county of Lincolnshire
13223|Cumbernauld||North Lanarkshire
13222||Notting Hill|the Royal Borough of Kensington and Chelsea
13217|Heigham||the city of Norwich
13216|Cheltenham||the county of Gloucestershire
13082|Home||
13081||Liverpool and of St James's|the city of Westminster
13080||Montgomery|the county of Powys and of Colomendy in the County of Clwyd
13079|Craighead||
13078|Breckland|Parson Cross|the county of South Yorkshire
13077|||
13076|Aberavon|Tandridge|the county of Surrey
13075|Idlicote|Shipston-on-Stow|the county of Warwickshire
13074|Guildford|Penton Mewsey|the county of Hampshire
13073|St Davids|Charlton|the London Borough of Greenwich
13349|Troon||the District of Kyle and Carrick
13350||Warrington|the county of Cheshire
13454|Woodside||the city of Aberdeen
13352|Chesterton||the county of Cambridgeshire
13353|Kings Heath|Birmingham|the county of West Midlands
13354|Tanworth|Stratford-upon-Avon|the county of Warwickshire
13355|Wirral||the county of Merseyside
13356|Westwell||the county of Oxfordshire
13341|North Bradley||the county of Wiltshire
13432|Lullington||the county of East Sussex
13486||Bresagh|the county of Down
13485|||
13488||New Romney|the county of Kent
13487||Richmond|the county of North Yorkshire
13490|||
13489|Lairg||the District of Sutherland
13339||Belgravia|the city of Westminster
13348|Holland Park|Southwold|the county of Suffolk
12963|Braunstone|Leicester|the county of Leicestershire
12859|Tullichettle|Comrie|the District of Perth and Kinross
12860|Paddington||the city of Westminster
12857||St Pancras|Greater London
12858|Jellicoe||
12863|Roding|Wanstead and Woodford|Greater London
12862||Liddington|the county of Wiltshire
10317||Deeside|the county of Clwyd
12866||Ainderby Quernhow|the county of North Yorkshire
12990||Bournville|the county of West Midlands
12989||Portsea|the county of Hampshire
12987||Ongar|the county of Essex
12994|The Shaws|Cathcart|the city of Glasgow
12993||Armagh|the county of Armagh
12992|Kincraig|Dysart|the District of Kirkcaldy
12991||Easton|the county of Leicestershire
10342|Bridgwater||the county of Somerset
13631|West Bromwich||the county of West Midlands
13634||Pemberton|the county of Lancashire
13218||Shrewsbury|the county of Shropshire
13219||Old Cantley|the county of South Yorkshire
13212||Kirkhill|the District of the city of Aberdeen
13213|Collingtree||the county of Northamptonshire
13214||Edgbaston|the county of West Midlands
13215|Dunphail||the District of Moray
13667||Artigarvan|the county of Tyrone
13668||Tewin|the county of Hertfordshire
13193|Lerwick||the Shetland Islands
13383|Horsell|Woking|the county of Surrey
13382|Monkton|Merrick and the Rhinns of Kells|Dumfries and Galloway
13377|Blaby|Newnham|the county of Northamptonshire
13376||Highgate|the London Borough of Haringey
13379|Crondall||the county of Hampshire
13378|Herne Hill||the London Borough of Southwark
13587|Portsoken||the city of London
13372||Mill Hill|the London Borough of Barnet
13649|Newnham||the county of Cambridgeshire
13647|Lindsay||
13648|Butterstone||
13645||Tooting|the London Borough of Wandsworth
13646|Listowel||
13297|Liverpool||
13298|Liverpool||
10365|Talgarth||the county of Powys
13296|Berwick|Ludlay|the county of East Sussex
13306|Highbury||the London Borough of Islington
13305||Sydmonton|the county of Hampshire
13132||Dewsbury|the county of West Yorkshire
13131|Pontefract||the county of West Yorkshire
13302|London||
13301|||
13300||Adur|the county of West Sussex
13299||Clerkenwell|the London Borough of Islington
13159|||
13154|||
12867|West Green||the county of Hampshire
12868|Bragar||the county of Ross and Cromarty
13562|||
13563||Churchhill|the District of the city of Edinburgh
13564|Dulwich|Bermondsey|the London Borough of Southwark
13565|Tradeston||the city of Glasgow
13566|Bearsden||the District of Bearsden and Milngavie
13567|Llandaff||the county of South Glamorgan
10386|Pulham Market||the county of Norfolk
12892|Haringey||Greater London
13121|Hudnall|Hampstead|the London Borough of Camden
13122|Clashfern|Eddrachillis|the District of Sutherland
13123|Drumadoon|Blackwaterfoot|the District of Cunninghame
13124|Culkein|Assynt|Highland
13125|Framwellgate|Durham|the county of Durham
13126|Benshie|Kirriemuir|the county of Angus
13127|Knebworth||the county of Hertfordshire
10396|Rogart||Sutherland
13129||Blackpool|the county of Lancashire
13130||Christchurch|the county of Dorset
10406|Drumglass|Carnteel|the county of Tyrone
12907||Studdridge|the county of Buckinghamshire
12905|||
12904|Mar||
12903|Mar and Kellie||Clackmannanshire
12902||Marlesford|the county of Suffolk
12901||Mannington|the county of Wiltshire
12910|Knightsbridge||the city of Westminster
12909|Ilton|Masham|the North Riding of the county of York
13551|Barnsley||South Yorkshire
13552|Darwen||the county of Lancashire
13549|Oxford||the county of Oxfordshire
13626|Twysden|Kilndown|the county of Kent
13632|||
10433|Gallanach|Oban|Argyll and Bute
13554|Chilthorne Domer||the county of Somerset
13546|Hendon|Gore|the London Borough of Barnet
13547||St Marylebone|the city of Westminster
13286||Hampstead|the London Borough of Camden
13285|Killead||the county of Antrim
13288|Langholm|Westerkirk|Dumfries and Galloway
13287|||
13290|Beaulieu||
13289|Montrose||
13276|Lower Marsh||the London Borough of Lambeth
13275|Wolvercote||the city of Oxford
13043|||
13044||Aberdyfi|the county of Gwynedd
13045|Huyton||the county of Merseyside
10446|Aberavon||the county of West Glamorgan and of Ceredigion in the County of Dyfed
13039|Manchester||the county of Greater Manchester
13040||Regents Park|the London Borough of Camden
13041|||
13042|||
13036|Lindisfarne|Hexham|the county of Northumberland
13705||Pateley Bridge|the county of North Yorkshire
13704||Sandy|the county of Bedfordshire
13703|Bladen|Briantspuddle|the county of Dorset
13702||Rothwell|the county of West Yorkshire
13709|Newcastle||
13708|Braintree|Coggeshall|the county of Essex
13689|Birkenhead||
13706|Winterbourne||the Royal county of Berkshire
13701||Renagour|the District of Stirling
13710||Newnham|the county of Cambridgeshire
13439||Goudhurst|the county of Sussex
13440||Brasted|the county of Kent
13438|||
13435|||
13436|Northesk||
13433||Telford|the county of Salop
13434||Cissbury|the county of West Sussex
13441|Louth||the county of Lincolnshire
13442|Seagrove Bay||the county of Isle of Wight
13165||The Barbican|the city of London
13164|Aylmerton||the county of Norfolk
13167|Bengarve|The Braid|the county of Antrim
13166|Onslow||
13161||Gloucester|the county of Gloucestershire
13163||Peckham Rye|the London Borough of Southwark
13162||the city of Plymouth|
13169||Liverpool|the county of Merseyside
13168|Oxford||
12945|||
12946||Walbrook|the city of London
12947||Kingston upon Hull|the East Riding of Yorkshire
12948|Monmouth|Broadway|the county of Hereford and Worcester
12949||Carnforth|the county of Lancashire
12951||Dunkeld|Perth and Kinross
12937|Blackburn|Langho|the county of Lancashire
12938||Wincanton|the county of Somerset
13603||Marylebone|the city of Westminster
13602|Rannoch|Bridge of Gaur|the District of Perth and Kinross
13601|||
10475||Stalybridge|the county of Greater Manchester
13009|Southwark|Charlbury|the county of Oxfordshire
13597||Mile End|Greater London
13596|Peterborough||
13595|Yeovil||the county of Somerset
13594|Sudbury||the county of Suffolk
12943|Worth Matravers|Belsize Park|the London Borough of Camden
13425|Oxenford|West Dowlish|the county of Somerset
13424||Caversham|the Royal county of Berkshire
13427|Highfield|Weelsby|the county of Humberside
13426|Writtle||the county of Essex
13429||Coleshill|the county of Warwickshire
13428|St Marylebone|the city of Westminster|
12916|Shulbrede||the county of West Sussex
12913|Portsmouth||
13695|Bayswater|Canterbury|the county of Kent
13071||Runnymede|the county of Surrey
13693||Brampton|the county of Suffolk
13694||Llanegryn|the county of Gwynedd
13699||Queensgate|the Royal Borough of Kensington and Chelsea
13700||Sandy|the county of Bedfordshire
13697||Holywell|the city of Oxford and county of Oxfordshire
13698||Bloomsbury|the London Borough of Camden
10495||Chester-le-Street|the county of Durham
13691|Cartvale||
13038|St Budeaux||the county of Devon
13037||Burnham Westgate|the county of Norfolk
13247|Ewell||the county of Surrey
13244||Mortlake|the London Borough of Richmond
13033|||
13032|||
13031||Redesdale|the county of Northumberland
13292||Goytre|the county of Gwent
13291||Hinton Blewitt|the county of Avon
12967|Babergh|Aldeburgh|the county of Suffolk
12970|Kaimsthorn|Hurlet|the District of Renfrew
13277||Wavertree|the county of Merseyside
13278||Huntingdon|the county of Cambridgeshire
13279|Mount Harry|Offham|the county of East Sussex
13280|Clifton|Chelsea|the Royal Borough of Kensington and Chelsea
13281||Ammanford|the county of Dyfed
13401|Calow||the county of Derbyshire
13405|Duntisbourne||the county of Gloucestershire
13332||Whitehall|the city of Westminster and of Hornsea in Yorkshire
13331|Conwy|Talyfan|the county of Gwynedd
10504|Port Ellen||
13333|Rochester||
13328|Earlsferry||the District of North East Fife
13327|Quarry Bank|Kentish Town|the London Borough of Camden
13330||Lower Iveagh|the county of Down
13329|Riverside|Chelsea|the Royal Borough of Kensington and Chelsea
10511||Perry Barr|the county of West Midlands
13005||Thorney Island|the city of Westminster
13006|Rosslyn||
13592|||
13590||Minginish|Highland
13588|Wensum||the county of Norfolk
13589||Staplefield|the county of West Sussex
13022|Preston Candover||the county of Hampshire
13026|Turville||the county of Buckinghamshire
12940|St Albans||
12939|St Edmundsbury and Ipswich||
13625|Bletso||
13624|Fawsley|Preston Capes|the county of Northamptonshire
13628|Salisbury||
12942|Abernethy||
12941||Passfield|the county of Hampshire
12912|Bowden|Melrose|the District of Ettrick and Lauderdale
13633|Sandwich||
13145|Newdigate||the county of Surrey
13146||Darlington|the county of Durham
13141|Asthal||the county of Oxfordshire
13142|Foscote||the county of Buckinghamshire
13143|Needham Market||the county of Suffolk
13144||Kineton|the county of Warwickshire
13181|Selborne||
13182|Douglas|Cramond|the city of Edinburgh
13184|||
13183||Gilcomstoun|the District of the city of Aberdeen
13186||Redlynch|the county of Wiltshire
13185|Guildford||the county of Surrey
13188||Chawton|Hampshire
13187|Northstead|Liversedge|the county of West Yorkshire
13189|Sheffield||
10535||Ashton-under-Lyne |the county of Greater Manchester
13191|Didgemere|Roydon|the county of Essex
13152|Shrewsbury||
13455|Greetland|Greetland and Stainland|the county of West Yorkshire
13456|||
13461|Glaisdale||the North Riding of the county of York
13462|Highbury|Canonbury|the London Borough of Islington
13459|Dunkeld||Perth and Kinross
13460|||
13463||Tilton|the county of East Sussex
13464|||
13653|Hadley|Eggington|the county of Bedfordshire
13654|Clifton|Mountsandel|the county of Londonderry
13324|Gilmorehill||the District of the city of Glasgow
13326|Leigh|Wigan|the county of Greater Manchester
13657|Snowdon||the county of West Sussex
13658|Swaffham Prior||the county of Cambridgeshire
13655|Southwark||
13656||St Pancras|the London Borough of Camden
13337|Aikwood|Ettrick Forest|The Scottish Borders
13338|Plaistow|Pall Mall|the city of Westminster
13385||Vauxhall|the London Borough of Lambeth
13384|Ludgate||the city of London
13387|Coddenham||the county of Suffolk
13386||Portmoak|the District of Perth and Kinross
13389||Swafield|the county of Norfolk
13557|Swindon|Reading|the Royal county of Berkshire
13627||Leyland|the county Palatine of Lancaster
13630|Blackheath||the London Borough of Greenwich
13629|||
13203|||
13204|Houndwood||the Scottish Borders
13205|||
13206|Vernham Dean||the county of Hampshire
13207||Tanlawhill|the county of Dumfries
13208||Pimlico|the city of Westminster
13209|Blackburn||the county of Lancashire
13194|Warwick||the county of Warwickshire
13195||Chingford|the London Borough of Waltham Forest
12978||White Lackington|the county of Somerset
10592||Llandaff|the county of South Glamorgan and of Leominster in the County of Herefordshire
12976|||
12975||Kesteven|the county of Lincolnshire
12974|Gresford||the county Borough of Wrexham
12973|Gwydir|Llanrwst|the county of Gwynedd
12972|Macclesfield|Prestbury|the county of Cheshire
12971|Swynnerton|Notting Hill|Greater London
12935|Walliswood|Dorking|the county of Surrey
12969|Monifieth||the District of the city of Dundee
13543||Manningham|the county of West Yorkshire
13544||Brailes|the county of Warwickshire
13541||Walsall|the county of West Midlands
13542||Sutton|the London Borough of Sutton
13539||Knutsford|the county of Cheshire
13540|||
13538||Sandwich|the county of Kent
13535|Truro||
13536||Widdington|the county of Essex
13272|||
13271|Camden||Greater London
13274||Bethnal Green|the London Borough of Tower Hamlets
13273|||
13268||Chesterfield|the county of Derbyshire
13267|Coleshill|Shrivenham|the county of Oxfordshire
13270||Roddam Dene|the county of Northumberland
13264||Read|the county of Lancashire
13263|Chorlton|Chester|the county of Cheshire
13114||Maldon|the county of Essex
13115|North Hill|Chewton Mendip|the county of Somerset
13117|Gestingthorpe||the county of Essex
13110|Worcester|Abbots Morton|the county of Hereford and Worcester
13112|Saltaire|Shipley|the county of West Yorkshire
13113||West Derby|the county of Merseyside
13119|||
13120|Detchant||the county of Northumberland
12896||Brockley|the London Borough of Lewisham
12895||Weeke|the city of Winchester
12894|Undercliffe||the county of West Yorkshire
12893|Invergowrie||Perth and Kinross
12900|Richmond||the London Borough of Richmond upon Thames
12899|||
12898||North East Croydon|the London Borough of Croydon
12897|Charlton|Highgate|Greater London
12888||Chelsea|Greater London
12957||Beeston|the county of Nottinghamshire
12958||Camberwell|the London Borough of Southwark
12961||Plymouth|the county of Devon
12962||Chesham Bois|the county of Buckinghamshire
12959|Crosby|Stevenage|the county of Hertfordshire
12960|Elvel|Llansantffraed|Elvel in the county of Powys
13617|Horton||the county of Somerset
13072|||
13616|Dinton||the county of Buckinghamshire
13619|Tillyorn|Finzean|the District of Kincardine and Deeside and of Fanling in Hong Kong
13618|Winchester||
13621||Windlesham|the county of Surrey
13620||Hammersmith|the London Borough of Hammersmith and Fulham
13623||Marylebone|the city of Westminster
13622|Sunningdale|Trevose|the county of Cornwall
13615||Barnes|the London Borough of Richmond
13614|Leeds||the county of West Yorkshire
12911|Worcester||
13025|Richmond|Richmond upon Thames|the London Borough of Richmond upon Thames
13023|Graffham||the county of West Sussex
13030|Old Scone||Perth and Kinross
13261|||
13293||Hampstead|the London Borough of Camden
13294||Kensington|the Royal Borough of Kensington and Chelsea
13197||Edgware|the London Borough of Barnet
13196||Moseley|the county of West Midlands
13548|Margravine|Barons Court|the London Borough of Hammersmith and Fulham
13545||Lancaster|the county of Lancashire
13201|Rising|Castle Rising|the county of Norfolk
13200|Chilton||the county of Suffolk
13199|Coles|Westmill|the county of Hertfordshire
13198|Bolton||the county of Greater Manchester
12845||St James's|the city of Westminster
13558|New Barnet||the London Borough of Barnet
13481||Ickenham|the London Borough of Hillingdon
13482||Aldgate|the city of London
13483||Southgate|the London Borough of Enfield
10554||Wednesbury|the county of West Midlands
13477|Llandudno||the county of Gwynedd
13478||Malone|the county of Antrim
13479||Oakley|Fife
13480|Drefelin||the county of Dyfed
13475||Battersea|the London Borough of Wandsworth
10425||Blackwaterfoot|Ayrshire and Arran
13055||Primrose Hill|the London Borough of Camden
13056||Mourne|the county of Down
13057|Luton||the county of Bedfordshire
13058||Mitcham and of Morden|the London Borough of Merton
13051||Harrow Weald|the London Borough of Harrow
13052||Fisherfield|Ross and Cromarty
13053|Brookwood||the county of Surrey
13054||Cambridge|the county of Cambridgeshire
13048|Hornsey||the London Borough of Haringey
10516||Merthyr Tydfil and of Rhymney|the county of Mid-Glamorgan
12838|Yarnbury||the county of Wiltshire
12837|Burry Port|Pembrey and Burry Port|the county of Dyfed
12836||Bracknell|the Royal county of Berkshire
12835||Rothiemay|Banffshire
12842||Killeen|the county of Down
12841|Eaton-under-Heywood||the county of Shropshire
12840|Richmond|Easby|the county of North Yorkshire
12839||Tottenham|the London Borough of Haringey
12844|Norwich||
12843|Tummel||Perth and Kinross
13449||Leeds|the county of West Yorkshire
13450|Norwood Green||the London Borough of Ealing
13447|Dillington||the county of Somerset
13448||Belfast|the county of Antrim
13445||Manchester|the county of Greater Manchester
13446||St Tudy|the county of Cornwall
13443|Kinlochard||Perth and Kinross
13444||Wychwood|the county of Oxfordshire
13452|Blaisdon||the county of Gloucestershire
13453|Leicester||
13175|Chelmsford||
13177|||
13176|Barnes||the London Borough of Richmond
13171||Bedwellty|the county of Gwent
13170|Glasgow||
13173|||
13172|||
13179|Thornes||the county of West Yorkshire
13178||Camden Town|the London Borough of Camden
13149||Kensington|the Royal Borough of Kensington and Chelsea
13150|Kirkwhelpington||the county of Northumberland
13151|Norfolk||
10345|Kirkhope||Scottish Borders
10584|Bolton||the county of Greater Manchester
10464|Clackmannan||Clackmannanshire
10612|||
10445|Yardley||the county of West Midlands
10291|Newport||the county of Gwent
10207|Bishop Auckland||the county of Durham
10101||Hamble-le-Rice|the county of Hampshire
10599||Kew|the London Borough of Richmond upon Thames
10211|Cumnock||East Ayrshire
10255|Epsom|West Anstey|the county of Devon
12928|Alamein||
10325|Cheltenham||the county of Gloucestershire
10536|Northwold||the county of Norfolk
10374|Markyate||the county of Hertfordshire
12933|Exeter||
13582||Bilston|the county of West Midlands
13583||Bennochy|Fife
10058|Nettlestone|St Helens|the county of Isle of Wight
10424||Peterborough|the county of Cambridgeshire
10110|Calton||the city of Edinburgh
10556||Hammersmith|the London Borough of Hammersmith and Fulham
10547|Finsbury||the London Borough of Islington
10003|Craigielea||Renfrewshire
13577||Gloucester|the county of Gloucestershire
10011|Swansea||the county of West Glamorgan
10135||St George|the county and city of Bristol
10234||Lincoln|the county of Lincolnshire
13319|Manchester||
10146|Felling||the county of Tyne and Wear
13321||Frognal|the London Borough of Camden
13320|Ecchinswell||the county of Hampshire
13323|Ludlow||the county of Shropshire
13322||Cumnor|the county of Oxfordshire
13315||Putney|the London Borough of Wandsworth
13714|York||
13174|Southwell and Nottingham||
13716||Enfield|the London Borough of Enfield
13718|Scarisbrick||the county of Lancashire
13717|Glen Clova||Angus
