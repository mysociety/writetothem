13375||Aldenham|the County of Shropshire
13368|||
13369||Thornes|the County of West Yorkshire
13370||Rotherham|the County of South Yorkshire
13371||Knock|the City of Belfast
13105|Megiddo||
13104||Norbury|the London Borough of Croydon
13103|Liverpool|Mossley Hill|the County of Merseyside
13102||Brondesbury|the London Borough of Brent
13109|||
13108||Southover|the County of East Sussex
13107|St Johns||the County of Surrey
13106|Sandwell||the County of West Midlands
13097|Weston-super-Mare||
13096|Ilminster|Ashill|the County of Somerset
12883|Arran||
12884||Chichester|the County of West Sussex
10015|Norton-sub-Hamdon||the County of Somerset
12882|Stoke|Widnes|the County of Cheshire
12879|Upholland|St Albans|the County of Hertfordshire
12880|||
12877|Hever||
12878||Richmond upon Thames|the London Borough of Richmond upon Thames
12875|||
12876|||
13526||Lutterworth|the County of Leicestershire
13525||Regent's Park|the City of Westminster
13528|Dorking|Iford|the County of East Sussex
13527|Bewdley||
13521|Tewkesbury|Gotherington|the County of Gloucestershire
13524||Anagach|Highland
13523||Heywood and Royton|Greater Manchester
13512|Brighton||the County of East Sussex
13503||Belgravia|the City of Westminster
13505||Cranford|the London Borough of Hilllingdon
13506|Craigweil||the County of West Sussex
13507||Godmanstone|the County of Dorset
13508||Hampton|the London Borough of Richmond
13510||Banbury|the County of Oxfordshire
13501|Cornhill|Boughrood|the County of Powys
13502||Liverpool|the County of Merseyside
13711|Crossharbour||the London Borough of Tower Hamlets
13241||Stoke Newington|Greater London
13240||Woodcote|the County of Surrey
13692||Blackwatertown|the County of Armagh
12981|Rowington||the County of Warwickshire
10054||Sandwell|the County of West Midlands
12980||Abbots Morton|the County of Hereford and Worcester
12985|Faversham||the County of Kent
12986||Warlingham|the County of Surrey and of Croydon in the London Borough of Croydon
12983||Pimlico|the City of Westminster
12984|Tara||
13028||Wallingford|the County of Oxfordshire
13034||Wigton|the County of Cumbria
13636||Bushfield|the County of Hampshire
13635||Bibury|the County of Gloucestershire
13638||Lydd|the County of Kent
13640|||
13639|||
13642||Lewes|the County of East Sussex
13610|Spennithorne||the County of North Yorkshire
13611|Alverthorpe||the County of West Yorkshire
10067|Sutton Mandeville||the County of Wiltshire
13613|||
13606||Ebbw Vale|the County of Gwent
13607|Tremorfa||the County of South Glamorgan
13608|||
13609|Madingley|Cambridge|the County of Cambridgeshire
13604||Camden|the London Borough of Camden
13430||Pitshanger|the London Borough of Ealing
13451||Goring|the County of Oxfordshire
13347|Brockwell|Herne Hill|the London Borough of Lambeth
13458||Rothley|the County of Leicestershire
13351|Caithness||
13676|Lochbroom||the District of Ross and Cromarty
13679|Alloway|Ayr|the District of Kyle and Carrick
10090||Allerdale|the County of Cumbria
13672|Canterbury||
13669|Clifton||the City and County of Bristol
13674|Berriew||the County of Powys
13670|Lour||the District of Angus
13018|Hadley|Monken Hadley|Greater London
13019||Upton|the County of Nottinghamshire
13017|Furness|Cartmel|the County of Cumbria
13014||Dean|the County of Oxfordshire
13015||Llantarnam|the County of Monmouth
13012|Wallasey|Leigh-on-Sea|the County of Essex
13010||Aldershot|the County of Hampshire
13253|Chester||
13252||Cranfield|the County of Bedfordshire
13251||Ryedale|the County of North Yorkshire
13258|Cholmondeley||
13257|||
13256||Leckhampton|the County of Gloucestershire
10108|Windermere||the County of Cumbria
13248|Hampstead||the London Borough of Camden
13517||Clapham|the London Borough of Lambeth
13518||Hackney|the London Borough of Hackney
13520|||
13514||Ranmore|the County of Surrey
13515|Pimlico||the City of Westminster
13516|Culross||
13550|||
13556||Langton Green|the County of Kent
12871|Berkeley||the County of Gloucestershire
10132|Castle Vale|Erdington|the County of West Midlands
12873|Courtown||
13235|Radley|Helhoughton|the County of Norfolk
13599|||
12952|||
12954|Crawford and Balcarres||
13094||Edgbaston|the County of West Midlands
13095||Pont Esgob|the Black Mountains and the County of Powys
13100||the London Borough of Croydon|
13098|Whitekirk||East Lothian
13099||Newick|the County of East Sussex
12966|Marylebone||the City of Westminster
13396|Coity|Penybont|the County of Mid Glamorgan
13395|Oldham|Broxbourne|the County of Hertfordshire
13393|Thornton-le-Fylde|Eccles|the County of Greater Manchester
13390|Alteryn||the County of Gwent
13659|||
13661||St Clement Danes|the City of Westminster
13662||Waltham Brooks|the County of West Sussex
13664||Jarrow|the County of Tyne and Wear
13665||Bocking|the County of Essex
13651||Ashton|the County of Northamptonshire
13000||Battersea|the London Borough of Wandsworth
12999|Dundee||
13002||Hong Kong Island|Hong Kong and of Knightsbridge in the Royal Borough of Kensington and Chelsea
12996|Durham||
12995||Armagh|the County of Armagh
12998||Stratton St Margaret|the County of Wiltshire
12997|Moulton||the County of North Yorkshire
13004|Winton|Rushyford|the County of Durham
13003||Kirkcaldy|Fife
13234||Nant Conwy|the County of Gwynedd
13232|Morpeth||the County of Northumberland and of the City of Newcastle upon Tyne
13233|||
13230||Aberteifi|the County of Dyfed
13231||Tunbridge Wells|the County of Kent and of Clerkenwell in the London Borough of Islington
13229|Erroll||
13242|Parkside|St Helens|the County of Merseyside
13243|Temple Guiting||the County of Gloucestershire
12852|Watford|Chipperfield|the County of Hertfordshire
12850||Horsham|the County of West Sussex
12851|Thoroton||the County of Nottinghamshire
12848||West Haddon|Northamptonshire
12849|||
12846|Ribbleton|Fulwood|the County of Lancashire
12847|Worcester|Wimbledon|the London Borough of Merton
10196||Southport|the County of Merseyside
12855||Frognal|the London Borough of Camden
13470||Shotesham|the County of Norfolk
13469|||
13472||Pimlico|the City of Westminster
13471|Llandaff||the County of South Glamorgan
13468|||
13467||Queen's Gate|the City of Westminster
13474||Plymouth|the County of Devon
13473|Drumlean||Stirling
13312|Thames Bank|Reddish|the County of Greater Manchester
10212||Sutton Coldfield|the County of West Midlands
13314|Carmyllie||the District of Angus
13307||Dingley|the County of Northamptonshire
13308|||
13309|Fairfield|Sauchie|the County of Clackmannanshire
13310||Blaenrhondda|the County of Mid Glamorgan
13304|Parkes|Southgate|Greater London and of Parkes in the State of New South Wales and Commonwealth of Australia
13063||Watford|the County of Hertfordshire
13062||Highgate|the London Borough of Camden
13061|||
13066|Market Rasen||the County of Lincolnshire
13065||Dudley|the County of West Midlands
13068||Glenridding|the County of Cumbria
12919|||
12920|||
12918|Chieveley||the Royal County of Berkshire
10233||Newcastle-under-Lyme|the County of Staffordshire
12924||Allerton|the County of Merseyside
12921||Youlbury|the County of Oxfordshire
12922|Strathblane|Deil's Craig|Stirling
12914|||
12915||Roundwood|the London Borough of Brent
13569|Potternewton|Leeds|the County of West Yorkshire
13568||Aldwych|the City of Westminster
13571|Edmonton||Greater London
13570|||
13572||Pendle|the County of Lancashire
13574||Ot Moor|the County of Oxfordshire
13561||Notting Hill|the Royal Borough of Kensington and Chelsea
13560|||
13415||Kilvey|the County of Swansea
13416||Govilon|the County of Gwent
13417|Fforestfach||the County of West Glamorgan
10247||Telford|the County of Shropshire
13420|Craigiebank||the City of Dundee
13421||Calverton|the County of Buckinghamshire
13422||Richmond upon Thames|the London Borough of Richmond upon Thames
13423||Kensington|the Royal Borough of Kensington and Chelsea
13140|Chiswick|Bedford Park|the London Borough of Ealing
13139||Chelmsford|the County of Essex
13137||Blackford|the City of Edinburgh
13135|Haringey|Hornsey|the London Borough of Haringey
13133|Peckham||the London Borough of Southwark
13148|Richmond||the County of North Yorkshire
13147||Chester|the County of Cheshire
13499||Higher Broughton|the County of Greater Manchester
13497||Sparkbrook|the County of West Midlands
13498||Isleworth|the London Borough of Hounslow
13495||Dartmouth Park|the London Borough of Camden
13496||Riddlesden|the County of West Yorkshire
13493|||
10276||Thenford|the County of Northamptonshire
13340||Worthing|the County of West Sussex
13224|Eggardon||the County of Dorset
13226|Astley Abbotts|Nash|the County of Shropshire
13221||Chedworth|the County of Gloucestershire
13220||Kettlethorpe|the County of Lincolnshire
13222||Notting Hill|the Royal Borough of Kensington and Chelsea
13217|Heigham||the City of Norwich
13082|Home||
13081||Liverpool and of St James's|the City of Westminster
13080||Montgomery|the County of Powys and of Colomendy in the County of Clwyd
13079|Craighead||
13078|Breckland|Parson Cross|the County of South Yorkshire
13077|||
13076|Aberavon|Tandridge|the County of Surrey
13075|Idlicote|Shipston-on-Stow|the County of Warwickshire
13074|Guildford|Penton Mewsey|the County of Hampshire
13073|St Davids|Charlton|the London Borough of Greenwich
13349|Troon||the District of Kyle and Carrick
13350||Warrington|the County of Cheshire
13454|Woodside||the City of Aberdeen
13352|Chesterton||the County of Cambridgeshire
13353|Kings Heath|Birmingham|the County of West Midlands
13355|Wirral||the County of Merseyside
13356|Westwell||the County of Oxfordshire
13432|Lullington||the County of East Sussex
13486||Bresagh|the County of Down
13485|||
13488||New Romney|the County of Kent
13487||Richmond|the County of North Yorkshire
13490|||
13489|Lairg||the District of Sutherland
13339||Belgravia|the City of Westminster
13348|Holland Park|Southwold|the County of Suffolk
12963|Braunstone|Leicester|the County of Leicestershire
12860|Paddington||the City of Westminster
12863|Roding|Wanstead and Woodford|Greater London
12862||Liddington|the County of Wiltshire
10317||Deeside|the County of Clwyd
12866||Ainderby Quernhow|the County of North Yorkshire
12990||Bournville|the County of West Midlands
12989||Portsea|the County of Hampshire
12994|The Shaws|Cathcart|the City of Glasgow
10589||Armagh|the County of Armagh
12992|Kincraig|Dysart|the District of Kirkcaldy
12991||Easton|the County of Leicestershire
10342|Bridgwater||the County of Somerset
13631|West Bromwich||the County of West Midlands
13634||Pemberton|the County of Lancashire
13219||Old Cantley|the County of South Yorkshire
13212||Kirkhill|the District of the City of Aberdeen
13213|Collingtree||the County of Northamptonshire
13214||Edgbaston|the County of West Midlands
13215|Dunphail||the District of Moray
13667||Artigarvan|the County of Tyrone
13668||Tewin|the County of Hertfordshire
13193|Lerwick||the Shetland Islands
13382|Monkton|Merrick and the Rhinns of Kells|Dumfries and Galloway
13377|Blaby|Newnham|the County of Northamptonshire
13376||Highgate|the London Borough of Haringey
13379|Crondall||the County of Hampshire
13378|Herne Hill||the London Borough of Southwark
13587|Portsoken||the City of London
13372||Mill Hill|the London Borough of Barnet
13649|Newnham||the County of Cambridgeshire
13647|Lindsay||
13648|Butterstone||
13645||Tooting|the London Borough of Wandsworth
13646|Listowel||
13297|Liverpool||
13298|Liverpool||
10365|Talgarth||the County of Powys
13296|Berwick|Ludlay|the County of East Sussex
13305||Sydmonton|the County of Hampshire
13132||Dewsbury|the County of West Yorkshire
13131|Pontefract||the County of West Yorkshire
13302|London||
13301|||
13300||Adur|the County of West Sussex
13299||Clerkenwell|the London Borough of Islington
13159|||
13154|||
12867|West Green||the County of Hampshire
12868|Bragar||the County of Ross and Cromarty
13562|||
13563||Churchhill|the District of the City of Edinburgh
13564|Dulwich|Bermondsey|the London Borough of Southwark
13565|Tradeston||the City of Glasgow
13566|Bearsden||the District of Bearsden and Milngavie
13567|Llandaff||the County of South Glamorgan
10386|Pulham Market||the County of Norfolk
12892|Haringey||Greater London
13121|Hudnall|Hampstead|the London Borough of Camden
13122|Clashfern|Eddrachillis|the District of Sutherland
13123|Drumadoon|Blackwaterfoot|the District of Cunninghame
13124|Culkein|Assynt|Highland
13125|Framwellgate|Durham|the County of Durham
13126|Benshie|Kirriemuir|the County of Angus
13127|Knebworth||the County of Hertfordshire
10396|Rogart||Sutherland
13129||Blackpool|the County of Lancashire
13130||Christchurch|the County of Dorset
10406|Drumglass|Carnteel|the County of Tyrone
12907||Studdridge|the County of Buckinghamshire
12905|||
12904|Mar||
12903|Mar and Kellie||Clackmannanshire
12902||Marlesford|the County of Suffolk
12901||Mannington|the County of Wiltshire
12910|Knightsbridge||the City of Westminster
12909|Ilton|Masham|the North Riding of the County of York
13551|Barnsley||South Yorkshire
13552|Darwen||the County of Lancashire
13549|Oxford||the County of Oxfordshire
13626|Twysden|Kilndown|the County of Kent
13632|||
13554|Chilthorne Domer||the County of Somerset
13546|Hendon|Gore|the London Borough of Barnet
13547||St Marylebone|the City of Westminster
13286||Hampstead|the London Borough of Camden
13285|Killead||the County of Antrim
13287|||
13290|Beaulieu||
13289|Montrose||
13276|Lower Marsh||the London Borough of Lambeth
13043|||
13044||Aberdyfi|the County of Gwynedd
13045|Huyton||the County of Merseyside
10446|Aberavon||the County of West Glamorgan and of Ceredigion in the County of Dyfed
13039|Manchester||the County of Greater Manchester
13040||Regents Park|the London Borough of Camden
13042|||
13705||Pateley Bridge|the County of North Yorkshire
13704||Sandy|the County of Bedfordshire
13703|Bladen|Briantspuddle|the County of Dorset
13702||Rothwell|the County of West Yorkshire
13709|Newcastle||
13708|Braintree|Coggeshall|the County of Essex
13689|Birkenhead||
13706|Winterbourne||the Royal County of Berkshire
13701||Renagour|the District of Stirling
13710||Newnham|the County of Cambridgeshire
13439||Goudhurst|the County of Sussex
13438|||
13435|||
13436|Northesk||
13433||Telford|the County of Salop
13434||Cissbury|the County of West Sussex
13441|Louth||the County of Lincolnshire
13442|Seagrove Bay||the County of Isle of Wight
13165||The Barbican|the City of London
13167|Bengarve|The Braid|the County of Antrim
13166|Onslow||
13161||Gloucester|the County of Gloucestershire
13163||Peckham Rye|the London Borough of Southwark
13162||the City of Plymouth|
13169||Liverpool|the County of Merseyside
12945|||
12946||Walbrook|the City of London
12947||Kingston upon Hull|the East Riding of Yorkshire
12949||Carnforth|the County of Lancashire
12951||Dunkeld|Perth and Kinross
12937|Blackburn|Langho|the County of Lancashire
12938||Wincanton|the County of Somerset
13603||Marylebone|the City of Westminster
13601|||
10475||Stalybridge|the County of Greater Manchester
13009|Southwark|Charlbury|the County of Oxfordshire
13597||Mile End|Greater London
13594|Sudbury||the County of Suffolk
12943|Worth Matravers|Belsize Park|the London Borough of Camden
13425|Oxenford|West Dowlish|the County of Somerset
13424||Caversham|the Royal County of Berkshire
13427|Highfield|Weelsby|the County of Humberside
13426|Writtle||the County of Essex
13429||Coleshill|the County of Warwickshire
12916|Shulbrede||the County of West Sussex
13695|Bayswater|Canterbury|the County of Kent
13071||Runnymede|the County of Surrey
13693||Brampton|the County of Suffolk
13694||Llanegryn|the County of Gwynedd
13699||Queensgate|the Royal Borough of Kensington and Chelsea
13697||Holywell|the City of Oxford and County of Oxfordshire
13698||Bloomsbury|the London Borough of Camden
10495||Chester-le-Street|the County of Durham
13691|Cartvale||
13038|St Budeaux||the County of Devon
13037||Burnham Westgate|the County of Norfolk
13244||Mortlake|the London Borough of Richmond
13033|||
13032|||
13031||Redesdale|the County of Northumberland
13291||Hinton Blewitt|the County of Avon
12967|Babergh|Aldeburgh|the County of Suffolk
12970|Kaimsthorn|Hurlet|the District of Renfrew
13277||Wavertree|the County of Merseyside
13279|Mount Harry|Offham|the County of East Sussex
13280|Clifton|Chelsea|the Royal Borough of Kensington and Chelsea
13281||Ammanford|the County of Dyfed
13401|Calow||the County of Derbyshire
13332||Whitehall|the City of Westminster and of Hornsea in Yorkshire
13331|Conwy|Talyfan|the County of Gwynedd
10504|Port Ellen||
13328|Earlsferry||the District of North East Fife
13327|Quarry Bank|Kentish Town|the London Borough of Camden
13330||Lower Iveagh|the County of Down
13329|Riverside|Chelsea|the Royal Borough of Kensington and Chelsea
10511||Perry Barr|the County of West Midlands
13005||Thorney Island|the City of Westminster
13006|Rosslyn||
13592|||
13588|Wensum||the County of Norfolk
13589||Staplefield|the County of West Sussex
13022|Preston Candover||the County of Hampshire
13026|Turville||the County of Buckinghamshire
13625|Bletso||
13624|Fawsley|Preston Capes|the County of Northamptonshire
13628|Salisbury||
12942|Abernethy||
12941||Passfield|the County of Hampshire
12912|Bowden|Melrose|the District of Ettrick and Lauderdale
13633|Sandwich||
13145|Newdigate||the County of Surrey
13146||Darlington|the County of Durham
13141|Asthal||the County of Oxfordshire
13142|Foscote||the County of Buckinghamshire
13143|Needham Market||the County of Suffolk
13144||Kineton|the County of Warwickshire
13181|Selborne||
13182|Douglas|Cramond|the City of Edinburgh
13184|||
13183||Gilcomstoun|the District of the City of Aberdeen
13186||Redlynch|the County of Wiltshire
13185|Guildford||the County of Surrey
13188||Chawton|Hampshire
13187|Northstead|Liversedge|the County of West Yorkshire
10535||Ashton-under-Lyne |the County of Greater Manchester
13191|Didgemere|Roydon|the County of Essex
13152|Shrewsbury||
13455|Greetland|Greetland and Stainland|the County of West Yorkshire
13456|||
13462|Highbury|Canonbury|the London Borough of Islington
13459|Dunkeld||Perth and Kinross
13460|||
13463||Tilton|the County of East Sussex
13464|||
13654|Clifton|Mountsandel|the County of Londonderry
13324|Gilmorehill||the District of the City of Glasgow
13326|Leigh|Wigan|the County of Greater Manchester
13657|Snowdon||the County of West Sussex
13658|Swaffham Prior||the County of Cambridgeshire
13337|Aikwood|Ettrick Forest|The Scottish Borders
13338|Plaistow|Pall Mall|the City of Westminster
13385||Vauxhall|the London Borough of Lambeth
13384|Ludgate||the City of London
13387|Coddenham||the County of Suffolk
13386||Portmoak|the District of Perth and Kinross
13389||Swafield|the County of Norfolk
13557|Swindon|Reading|the Royal County of Berkshire
13630|Blackheath||the London Borough of Greenwich
13629|||
13203|||
13204|Houndwood||the Scottish Borders
13205|||
13206|Vernham Dean||the County of Hampshire
13207||Tanlawhill|the County of Dumfries
13208||Pimlico|the City of Westminster
13209|Blackburn||the County of Lancashire
13194|Warwick||the County of Warwickshire
13195||Chingford|the London Borough of Waltham Forest
12978||White Lackington|the County of Somerset
10592||Llandaff|the County of South Glamorgan and of Leominster in the County of Herefordshire
12976|||
12975||Kesteven|the County of Lincolnshire
12974|Gresford||the County Borough of Wrexham
12972|Macclesfield|Prestbury|the County of Cheshire
12971|Swynnerton|Notting Hill|Greater London
12935|Walliswood|Dorking|the County of Surrey
13543||Manningham|the County of West Yorkshire
13544||Brailes|the County of Warwickshire
13541||Walsall|the County of West Midlands
13542||Sutton|the London Borough of Sutton
13539||Knutsford|the County of Cheshire
13540|||
13538||Sandwich|the County of Kent
13536||Widdington|the County of Essex
13272|||
13271|Camden||Greater London
13274||Bethnal Green|the London Borough of Tower Hamlets
13273|||
13267|Coleshill|Shrivenham|the County of Oxfordshire
13270||Roddam Dene|the County of Northumberland
13264||Read|the County of Lancashire
13263|Chorlton|Chester|the County of Cheshire
13114||Maldon|the County of Essex
13115|North Hill|Chewton Mendip|the County of Somerset
13117|Gestingthorpe||the County of Essex
13110|Worcester|Abbots Morton|the County of Hereford and Worcester
13112|Saltaire|Shipley|the County of West Yorkshire
13113||West Derby|the County of Merseyside
13119|||
13120|Detchant||the County of Northumberland
12896||Brockley|the London Borough of Lewisham
12895||Weeke|the City of Winchester
12894|Undercliffe||the County of West Yorkshire
12893|Invergowrie||Perth and Kinross
12900|Richmond||the London Borough of Richmond upon Thames
12899|||
12888||Chelsea|Greater London
12957||Beeston|the County of Nottinghamshire
12958||Camberwell|the London Borough of Southwark
12961||Plymouth|the County of Devon
12962||Chesham Bois|the County of Buckinghamshire
12959|Crosby|Stevenage|the County of Hertfordshire
12960|Elvel|Llansantffraed|Elvel in the County of Powys
13617|Horton||the County of Somerset
13616|Dinton||the County of Buckinghamshire
13619|Tillyorn|Finzean|the District of Kincardine and Deeside and of Fanling in Hong Kong
13618|Winchester||
13621||Windlesham|the County of Surrey
13620||Hammersmith|the London Borough of Hammersmith and Fulham
13623||Marylebone|the City of Westminster
13622|Sunningdale|Trevose|the County of Cornwall
13615||Barnes|the London Borough of Richmond
13614|Leeds||the County of West Yorkshire
13025|Richmond|Richmond upon Thames|the London Borough of Richmond upon Thames
13023|Graffham||the County of West Sussex
13030|Old Scone||Perth and Kinross
13294||Kensington|the Royal Borough of Kensington and Chelsea
13197||Edgware|the London Borough of Barnet
13196||Moseley|the County of West Midlands
13548|Margravine|Barons Court|the London Borough of Hammersmith and Fulham
13545||Lancaster|the County of Lancashire
13201|Rising|Castle Rising|the County of Norfolk
13200|Chilton||the County of Suffolk
13199|Coles|Westmill|the County of Hertfordshire
13198|Bolton||the County of Greater Manchester
12845||St James's|the City of Westminster
13558|New Barnet||the London Borough of Barnet
13481||Ickenham|the London Borough of Hillingdon
13482||Aldgate|the City of London
13483||Southgate|the London Borough of Enfield
10554||Wednesbury|the County of West Midlands
13477|Llandudno||the County of Gwynedd
13478||Malone|the County of Antrim
13479||Oakley|Fife
13480|Drefelin||the County of Dyfed
13475||Battersea|the London Borough of Wandsworth
10425||Blackwaterfoot|Ayrshire and Arran
13055||Primrose Hill|the London Borough of Camden
13056||Mourne|the County of Down
13057|Luton||the County of Bedfordshire
13058||Mitcham and of Morden|the London Borough of Merton
13051||Harrow Weald|the London Borough of Harrow
13052||Fisherfield|Ross and Cromarty
13053|Brookwood||the County of Surrey
13054||Cambridge|the County of Cambridgeshire
13048|Hornsey||the London Borough of Haringey
10516||Merthyr Tydfil and of Rhymney|the County of Mid-Glamorgan
12838|Yarnbury||the County of Wiltshire
12837|Burry Port|Pembrey and Burry Port|the County of Dyfed
12836||Bracknell|the Royal County of Berkshire
12835||Rothiemay|Banffshire
12842||Killeen|the County of Down
12841|Eaton-under-Heywood||the County of Shropshire
12840|Richmond|Easby|the County of North Yorkshire
12839||Tottenham|the London Borough of Haringey
12844|Norwich||
12843|Tummel||Perth and Kinross
13450|Norwood Green||the London Borough of Ealing
13447|Dillington||the County of Somerset
13445||Manchester|the County of Greater Manchester
13443|Kinlochard||Perth and Kinross
13444||Wychwood|the County of Oxfordshire
13452|Blaisdon||the County of Gloucestershire
13453|Leicester||
13177|||
13176|Barnes||the London Borough of Richmond
13171||Bedwellty|the County of Gwent
13170|Glasgow||
13173|||
13172|||
13179|Thornes||the County of West Yorkshire
13178||Camden Town|the London Borough of Camden
13149||Kensington|the Royal Borough of Kensington and Chelsea
13150|Kirkwhelpington||the County of Northumberland
13151|Norfolk||
10345|Kirkhope||Scottish Borders
10584|Bolton||the County of Greater Manchester
10464|Clackmannan||Clackmannanshire
10612|||
10445|Yardley||the County of West Midlands
10291|Newport||the County of Gwent
10207|Bishop Auckland||the County of Durham
10101||Hamble-le-Rice|the County of Hampshire
10599||Kew|the London Borough of Richmond upon Thames
10211|Cumnock||East Ayrshire
10255|Epsom|West Anstey|the County of Devon
12928|Alamein||
10325|Cheltenham||the County of Gloucestershire
10536|Northwold||the County of Norfolk
10374|Markyate||the County of Hertfordshire
12933|Exeter||
10607||Bilston|the County of West Midlands
13583||Bennochy|Fife
10058|Nettlestone|St Helens|the County of Isle of Wight
10424||Peterborough|the County of Cambridgeshire
10110|Calton||the City of Edinburgh
10556||Hammersmith|the London Borough of Hammersmith and Fulham
10547|Finsbury||the London Borough of Islington
10003|Craigielea||Renfrewshire
13577||Gloucester|the County of Gloucestershire
10011|Swansea||the County of West Glamorgan
10135||St George|the County and City of Bristol
10234||Lincoln|the County of Lincolnshire
13682|Manchester||
10146|Felling||the County of Tyne and Wear
13321||Frognal|the London Borough of Camden
13320|Ecchinswell||the County of Hampshire
13323|Ludlow||the County of Shropshire
13322||Cumnor|the County of Oxfordshire
13315||Putney|the London Borough of Wandsworth
13714|York||
13716||Enfield|the London Borough of Enfield
13718|Scarisbrick||the County of Lancashire
13717|Glen Clova||Angus
13500||Skidby|the County of the East Riding of Yorkshire
10136||Congresbury|the County of Somerset
13720|Holbeach|South Holland|the County of Lincolnshire
13721||Whitcurch|the County of Devon
13724|Trafford|Bowdon|the County of Cheshire
13723||Odstock|the County of Wiltshire
13725||Gateshead|the County of Tyne and Wear
13727|Handsworth|Handsworth|the County of West Midlands
13728|Winchester|Winchester|the County of Hampshire
13726||Holland Park|the Royal Borough of Kensington and Chelsea
13730||Leicester|the County of Leicestershire
13729|Fairford|Fairford|the County of Gloucestershire
13731||Eaglescliffe|the County of Durham
13732||Tregony|the County of Cornwall
13734||Cornhill|the City of London
13733||Clogher Valley|the County of Tyrone
13737|St George's||the County of Antrim
13740||Cunninghame|North Ayrshire
13739|Bradford||the County of West Yorkshire
13876|Dalston||the London Borough of Hackney
13877|Whitchurch||the County of South Glamorgan
10059||Withington|the County of Greater Manchester
13880|Blackheath|Wild Brooks|the County of West Sussex
13882||Kilgetty|the County of Dyfed
13878|Belmont|Belmont|the County of Antrim
13881||Chelsea|the Royal Borough of Kensington and Chelsea
13879||Marsh Green|the County of Devon
13168|Pentregarth|Ceinewydd|the County of Dyfed
13883|Ripon and Leeds||
13884||Willersey|the County of Gloucestershire
13885||Spitalfields|the London Borough of Tower Hamlets
13886|Ewelme|Ewelme|the County of Oxfordshire
12897|Charlton|Highgate|Greater London
13738|Duncansby||Caithness
13602|Rannoch|Bridge of Gaur|the District of Perth and Kinross
13072|||
13890|Aldringham||the County of Suffolk
13920|Abbotsbury||the County of Dorset
13919|||
13922||Whitehall Park|the London Borough of Islington
13921|Surbiton||the Royal Borough of Kingston-upon-Thames
13923||Hampstead|the London Borough of Camden
13924||Wytham|the County of Oxfordshire
13925||Bromley-by-Bow|the London Borough of Tower Hamlets
13926||Donegore|the County of Antrim
13929||St Leonard's Forest|the County of West Sussex
13928|Spithead|Seaview|the County of Isle of Wight
13931||Holland Park|the Royal Borough of Kensington and Chelsea
13559||Queensbury|Greater London
13932|Denham|Gerrards Cross|the County of Buckinghamshire
13937||Dewsbury|the County of West Yorkshire
13936||Hutton Roof|the County of Cumbria
13939||Chalford Hill|the County of Gloucestershire
13938|Frognal|Hampstead|the London Borough Camden
13940|Tankerness||Orkney
10605||Lisnagarvey|the County of Antrim
14126||Heslington|the County of North Yorkshire
14125|Brentford|Elsted|the County of West Sussex and of Wimbledon in the London Borough of Merton
14127|Chichester||
14129|Stair||
14130||Queen's Park|the County of East Sussex
14132|Lincoln||
14133||Northampton|the County of Northamptonshire
14134||Langbaurgh|the County of North Yorkshire
14135|Bath and Wells||
13261|Salisbury||
14136|Kelvin||the City of Glasgow
14138||Draycote|the County of Warwickshire
10412||Foy|the County of Herefordshire and of Hartlepool in the County of Durham
14139|Barnes||the London Borough of Richmond upon Thames
14140||Truro|the County of Cornwall
14143||Radlett|the County of Hertfordshire
14144|Bradford||
14145|Abersoch||the County of Gwynedd
14147|Loughborough||the County of Leicestershire
24686|Mapesbury|Hampstead Town|the London Borough of Camden
24685|Stone-cum-Ebony||the County of Kent
24687|Wakefield||
24688|Tonaghmore||the County of Down
24689||Eastry|the County of Kent
13930|Birmingham|Alvechurch and of Bromsgrove|the County of Worcestershire
24690|Holyhead||the County of Ynys M�n
24693|Bristol||
24692||Clapton|the London Borough of Hackney
10420|Springburn|Port Dundas|the City of Glasgow
24694||Kirkinriola|the County of Antrimsgow
24695||Aldgate|the City of London
24696|||
24700|Blackburn||
24699|Lichfield||
24698|Hereford||
24706|Gloucester||
24705|Birkenhead||the County of Cheshire
24704||Loxbeare|the County of Devon
