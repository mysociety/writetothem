13375|30 July 1941|Trinity College, Oxford
13368|24 August 1963|Aberdeen University
13369|21 July 1962|Polytechnic of East London
13370|24 April 1957|Thomas Rotherham College, Rotherham; Sheffield Hallam University
13371|28 March 1955|Queen's University, Belfast
13105|20 April 1931|RMA, Sandhurst
13104|16 November 1964|
13103|15 March 1951|Christ's College, Liverpool; St Andrews University
13102|13 March 1954|Warwick University; Birmingham University; University of East Anglia
13109|15 October 1921|
13108|16 May 1943|University College of Wales, Aberystwyth; Sussex University
13107|17 July 1947|Bristol University; London University Institute of Education; Brunel University
13106|20 November 1926|London School of Economics; University College, London
13097|15 April 1940|Brasenose College, Oxford
13096|30 March 1927|Christ Church, Oxford
12883|14 July 1938|Balliol College, Oxford
12884|4 March 1946|
10015|27 February 1941|
12882|6 December 1922|Ruskin College, Oxford; Gonville and Caius College, Cambridge
12879|20 March 1956|Bedford College, London University
12880|27 December 1951|
12877|16 June 1946|
12878|29 August 1923|Leverhulme scholarship to Royal Academy of Dramatic Art
12875|3 October 1956|
12876|29 September 1928|Balliol College, Oxford
13526|25 December 1946|New College, Oxford
13525|24 August 1930|
13528|3 November 1934|Magdalen College, Oxford
13527|3 January 1938|Trinity College, Cambridge
13521|17 June 1918|Royal Agricultural College, Cirencester
13524|31 January 1961|Southampton University
13523|14 October 1923|Correspondence course, qualified as Accountant
13512|11 June 1953|Sussex University; Kent University
13503|18 October 1941|
13505|20 September 1939|Trinity College, Cambridge
13506|15 March 1936|St John's College, Cambridge
13507|22 June 1945|Nottingham University
13508|18 March 1932|
13510|31 July 1939|College of Education (London); Department of Education, Oxford University
13501|13 October 1933|Balliol College, Oxford
13502|10 December 1944|St Catherine's College, Oxford
13711|25 August 1944|Carleton University, Canada; Laval University, Canada; McGill University, Canada
13241|27 September 1942|London School of Economics
13240|29 July 1952|Trinity College, Cambridge; Wharton Business School, University of Pennsylvania
13692|26 May 1938|
12981|8 May 1940|Glasgow University
10054|8 October 1929|Dewsbury College of Commerce and Art
12980|13 March 1931|Manchester University
12985|21 March 1930|King's College, London University
12986|19 May 1943|Law Society School of Law, College of Law
12983|2 April 1943|Britannia Royal Naval College, Dartmouth
12984|20 December 1946|
13028|9 September 1936|Reading University
13034|6 October 1939|Wadham College, Oxford
13636|18 December 1923|Army Staff College; Imperial Defence College
13635|19 March 1942|Manchester University
13638|6 March 1942|
13640|5 December 1930|
13639|27 November 1927|New College, Oxford
13642|7 May 1921|Sidney Sussex College, Cambridge; London School of Economics
13610|25 September 1939|Trinity College, Cambridge; Yale University, USA
13611|21 June 1942|
10067|3 March 1934|Balliol College, Oxford; Harvard Business School; Commonwealth (Harkness) Fund Fellow, Harvard
13613|30 June 1952|Royal Agricultural College, Cirencester
13606|3 January 1937|
13607|12 April 1927|Coleg Harlech
13608|2 August 1938|Northampton Institute of Agriculture
13609|20 February 1948|St John's College, Cambridge; Stanford University, USA
13604|30 March 1930|Magdalen College, Oxford
13430|13 March 1944|Manchester University
13451|12 March 1954|Inns of Court School of Law; Columbia Law School, New York
13347|3 January 1938|University College, Oxford
13458|14 January 1941|Moulton Agricultural College, Northampton
13351|3 November 1948|Royal Agricultural College, Cirencester
13676|11 June 1931|Corpus Christi, Oxford; Edinburgh University
13679|24 May 1917|Ecole des Sciences Politiques, Paris 1934; Trinity Hall, Cambridge
10090|23 August 1943|The Sorbonne, Paris
13672|14 June 1950|Christ's College, Cambridge; Christ Church and Wadham Colleges, Oxford
13669|13 November 1935|King's College, London; London College of Divinity
13674|12 February 1948|King's College, London University; Council of Legal Education
13670|28 April 1925|
13018|11 November 1916|Gonville and Caius College, Cambridge
13019|6 June 1919|RMC, Sandhurst
13017|2 November 1941|
13014|24 August 1942|Selwyn College, Cambridge
13015|5 December 1919|School of Slavonic Studies, London University
13012|29 April 1942|Heidelberg University; London University; Central London Polytechnic
13010|12 February 1953|Worcester College, Oxford
13253|16 March 1950|Merton College, Oxford; Edinburgh University
13252|30 October 1926|Bristol University
13251|1 May 1936|Birmingham University; University of Kansas
13258|27 June 1960|Sorbonne
13257|14 August 1930|Gonville and Caius College, Cambridge
13256|25 April 1925|Westminster College of Commerce
10108|19 October 1939|Manchester University; Sheffield University
13248|17 April 1932|Ruskin College, Oxford
13517|26 October 1949|Trinity College, Cambridge
13518|6 December 1928|King's College, London University
13520|14 July 1937|Trinity College, Cambridge
13514|29 September 1956|Loughborough University
13515|4 July 1940|Newnham College, Cambridge
13516|19 July 1933|New College, Oxford
13550|1 January 1942|St Bartholomew's Hospital and Royal Dental Hospital, London University
13556|10 March 1947|St Peter's College, Oxford
12871|13 May 1937|
10132|22 December 1933|
12873|19 March 1954|Berkshire College of Agriculture; Royal Agricultural College, Cirencester
13559|6 July 1937|London Hospital; London University external student
13235|17 September 1929|Lincoln College, Oxford
13599|9 June 1944|London University
12952|12 September 1939|Trinity College, Cambridge
12954|5 March 1927|Trinity College, Cambridge
13094|9 January 1950|Digby Stuart Training College, Roehampton
13095|25 February 1934|Trinity College, Cambridge
13100|15 December 1917|London School of Economics statistics 1938
13098|18 November 1935|St Andrews University; Edinburgh University
13099|27 January 1943|
12966|9 December 1946|Manchester University; Birmingham University; London University
13396|24 June 1935|Bridgend Technical College
13395|9 November 1939|University College, London; Institute of Education; London School of Economics
13393|29 April 1943|
13390||
13659|3 October 1927|King's College, Cambridge
13661|10 July 1940|University of Bombay; University of Pennsylvania
13662|4 March 1937|Institute of Science, Bhavnager, Gujarat, India; Brighton Technical College
13664|6 March 1929|
13665|30 September 1934|Writtle Agricultural College, Essex
13651|8 September 1934|Lincoln College, Oxford; Nuffield College, Oxford; Harvard University, USA
13000|5 December 1932|London School of Economics
12999|5 June 1949|St Andrews University
13002|29 February 1940|College of the Holy Names, Oakland, California; University of California, Berkeley, California
12996|1 December 1948|Exeter College, Oxford
12995|27 April 1937|Queen's University, Belfast; Trinity College, Dublin
12998|2 February 1945|Queens' College, Cambridge; Harvard University
12997|4 October 1933|Open University
13004|15 September 1925|
13003|9 May 1950|Edinburgh University
13234|18 October 1946|University College of Wales
13232|11 December 1920|
13233|2 March 1930|New College, Oxford
13230|7 December 1932|University of Wales, Aberystwyth
13231|10 September 1935|St George's Hospital; Battersea College of Technology
13229|20 April 1948|Trinity College, Cambridge
13242|19 October 1930|
13243|7 August 1941|London School of Economics
12852|30 November 1942|Watford College of Technology
12850|23 February 1919|Magdalene College, Cambridge
12851|19 November 1951|Queens' College, Cambridge
12848|10 March 1932|Queen Mary College, London University
12849|8 May 1935|
12846|29 June 1940|
12847|22 March 1946|Worcester College, Oxford
10196|6 February 1931|
12855|23 September 1926|SE London Technical College
13470|11 December 1941|
13469|8 June 1929|Magdalene College, Cambridge
13472|1 July 1944|Clare College, Cambridge; Manchester University; Birmingham University
13471|23 February 1949|St Mary's Hospital, London University
13468|13 February 1934|University College, London
13467|13 September 1924|Gonville and Caius College, Cambridge; Birmingham University
13474|21 February 1936|Royal Holloway College, London University
13473|16 October 1954|St Andrews University
13312|1 June 1935|School of Architecture, Manchester University; School of Architecture, Yale University; Henry Fellowship and Guest Fellow, Jonathan Edwards College, Yale School of Architecture 1962
10212|2 February 1938|Trinity Hall, Cambridge
13314|29 May 1945|Gonville and Caius College, Cambridge; Edinburgh University
13307|27 May 1942|Balliol College, Oxford; Institute of Chartered Accountants, England and Wales
13308|15 December 1970|Camberwell College of Arts 1989-94
13309|10 April 1941|Co-operative College, Loughborough
13310|28 November 1940|Pontypridd Technical College 1970-73; University College of Wales, Cardiff
13304|17 July 1927|East Sydney Technical College; Sydney University; Cordon Bleu de Paris
13063|28 February 1941|Madrid University
13062|13 September 1930|St Peter's College, Oxford
13061|3 September 1937|Gonville and Caius College, Cambridge; Harvard Business School 1969
13066|10 December 1940|Chelmsford College of Further Education; Essex University
13065|5 April 1927|St John's College, Oxford; New York University
13068|17 December 1912|Bede College, Durham
12919|7 October 1944|
12920|21 April 1935|Grenoble University, France
12918|12 November 1926|New College, Oxford
10233|21 March 1933|Cardiff Royal Infirmary School of Radiography
12924|5 January 1950|Gonville and Caius College, Cambridge; University College, London
12921|18 January 1933|Trinity College, Cambridge; Harvard Law School
12922|17 May 1936|Glasgow University
12914|16 November 1965|
12915|2 September 1946|
13569|29 October 1932|Bradford Technical College
13568|21 March 1945|London School of Economics; Lincoln's Inn
13571|26 March 1925|WEA Co-operative College 1964; Open University
13570|8 April 1951|London School of Economics
13572|27 July 1942|Hertford College, Oxford
13574|1 October 1950|St Hilda's College, Oxford; Honorary Fellowship, St Hilda's College, Oxford 1999
13561|29 June 1935|London School of Economics
13560|21 May 1941|
13415|23 May 1935|King's College, Cambridge 1959
13416|26 September 1923|St John's College, Cambridge
13417|27 December 1941|London School of Economics
10247|1 November 1940|Leicester University; Manchester University
13420|17 November 1938|Royal Military Academy, Sandhurst
13421|23 June 1927|King's College, Cambridge; Cuddesdon Theological College, Oxford
13422|12 January 1947|Girton College, Cambridge
13423|23 September 1939|
13140|28 September 1935|New College, Oxford
13139|16 September 1940|Nuffield Scholarship for Agriculture
13137|8 January 1946|Edinburgh University
13135|11 October 1953|Trinity College, Cambridge
13133|15 September 1942|
13148|4 January 1944|Ealing Hotel and Catering College
13147|28 September 1947|Warwick University; Sussex University; Keele University
13499|8 October 1934|Salford College of Advanced Technology
13500|30 May 1937|Trinity College, Dublin
13497|28 December 1932|Hull University
13498|8 August 1925|Croydon and Borough Polytechnics
13495|26 March 1949|Newnham College, Cambridge
13496|30 August 1917|Balliol College, Oxford
13493|22 November 1953|Durham University
10276|21 March 1933|Pembroke College, Oxford
13340|18 January 1928|Gonville and Caius College, Cambridge; Yale University, USA
13224|12 January 1936|Manchester University 1971; London University
13226|25 April 1942|Oxford University; Wharton School of Finance, Pennsylvania University
13221|8 May 1934|University of Cape Town; The Queen's College, Oxford
13220|14 May 1946|Lady Margaret Hall, Oxford
13222|20 May 1945|Nottingham University
13217|24 May 1941|Cambridge University; University of California and Columbia University, New York; Nuffield College, Oxford
13082|20 November 1943|Christ Church, Oxford
13081|25 May 1939|Royal Ballet School; Southampton University; Universidad Central, Ecuador
13080|26 March 1925|University College of Wales, Aberystwyth; Gray's Inn
13079|27 June 1938|St John's College, Cambridge; Edinburgh University
13078|5 September 1940|Leicester University
13077|29 January 1951|Christ Church, Oxford
13076|20 December 1926|Trinity Hall, Cambridge
13075|8 February 1932|London School of Economics
13074|18 January 1936|King's College, Cambridge
13073|10 Jan 1931|
13349|2 March 1924|Royal Technical College, Glasgow
13350|17 February 1930|Horwich Technical College
13454|3 January 1932|
13352|5 September 1941|Trinity College, Cambridge; Warwick University
13353|19 May 1949|Leeds University
13355|21 May 1942|Montpellier University, France; Bristol University; Guildford College of Law
13356|8 March 1930|Trinity College, Cambridge
13432|28 March 1915|Magdalen College, Oxford
13486|29 June 1931|Balliol College, Oxford; Queen's University, Belfast
13485|13 June 1932|Trinity College, Oxford
13488|27 April 1933|Holborn College of Law, Languages and Commerce
13487|5 August 1935|RMA, Sandhurst
13490|31 July 1951|Trinity College, Cambridge; Cumbria College of Agriculture and Forestry
13489|23 June 1940|Glasgow University; Christ's College, Cambridge
13339|13 November 1931|London University
13348|3 August 1920|
12963|11 July 1928|Trinity Hall, Cambridge; Harvard Post-Graduate Law School, USA 1953
12860|18 November 1939|Somerville College, Oxford
12863|7 September 1926|Jesus College, Cambridge
12862|12 May 1932|University of Witwatersrand
10317|26 June 1937|Teacher training, Normal College, Bangor, North Wales
12866|10 December 1930|King's College, Newcastle upon Tyne
12990|28 January 1936|
12989|28 March 1935|London School of Economics
12994|12 May 1950|Council of Legal Education
10589|24 December 1937|Queen's University, Belfast
12992|29 July 1926|Edinburgh University
12991|18 October 1928|Trinity College, Cambridge
10342|13 June 1933|Emmanuel College, Cambridge
13631|24 April 1937|Punjab University, India; National Foundry College, Wolverhampton; Aston University, Birmingham; Teacher Training College, Wolverhampton; Essex University
13634|5 January 1927|Trinity College, Oxford
13219|14 December 1944|
13212|7 May 1930|
13213|9 July 1927|
13214|3 October 1920|Police Staff College
13215|12 May 1923|Jesus College, Cambridge
13667|23 April 1944|
13668|19 July 1936|Durham University; Rainer House 1960-61; London School of Economics 1964-65
13193|8 May 1942|Fitzwilliam College, Cambridge
13382|27 June 1940|Sidney Sussex College, Cambridge
13377|11 March 1932|Christ Church, Oxford
13376|15 March 1934|King's College, Cambridge; London School of Economics
13379|2 November 1937|Christ's College, Cambridge
13378|3 July 1936|Trinity College, Cambridge; Harvard Law School
13587|8 December 1941|Manchester University
13372|11 July 1944|F.C.A. 1966
13649|13 February 1928|London University; Nottingham University; Manchester University; Sidney Sussex College, Cambridge
13647|19 November 1955|Edinburgh University; University of California, Davis
13648|15 April 1943|Sussex University; London University
13645|21 April 1948|Magdalen College, Oxford
13646|28 June 1964|Queen Mary and Westfield College, London
13297|18 August 1948|Exeter University; PGCE in drama and RE 1971; Wycliffe Hall, Oxford 1982
13298|14 November 1944|Perugia University, Italy
10365|2 May 1935|Seale Hayne Agricultural College; Reading University
13296|9 May 1929|Trinity College, Cambridge; Harvard Law School
13305|22 March 1948|Magdalen College, Oxford; Royal College of Music
13132|22 January 1924|Ruskin College, Oxford
13131|18 December 1925|Leeds University
13302|11 July 1947|Trinity College, Cambridge; Cuddesdon Theological College, Oxford; Lincoln Theological College
13301|7 Jun 1951|
13300|14 October 1936|Christ's College, Cambridge; Wadham College, Oxford
13299|14 March 1951|London School of Economics: international history 1972,  European studies; Inns of Court School of Law
13159|13 January 1933|Trinity College, Cambridge
13154|27 March 1939|Christ Church, Oxford
12867|14 May 1942|
12868|14 November 1933|Glasgow University
13562|30 July 1925|Ruskin College, Oxford; Merton College, Oxford; Nuffield College, Oxford
13563|12 June 1929|Edinburgh University
13564|6 January 1933|London University
13565|20 August 1940|l.c.m Apprenticeship, marine engineer
13566|5 March 1926|
13567|1 April 1926|Bedford and Birkbeck Colleges, London University 1967, HV Tut Cert 1960
10386|14 February 1937|St Andrews University; King's College, London University
12892|30 April 1933|Jesus College, Oxford; Ohio State University
13121|23 September 1946|York University
13122|2 July 1927|Edinburgh University; Trinity College, Cambridge
13123|30 January 1946|Edinburgh University; University of Virginia, USA
13124|25 February 1940|Leverndale School of Nursing, Glasgow; West Cumberland School of Nursing, Whitehaven
13125|21 March 1943|London University; FBI National Academy, Quantico, USA
13126|10 July 1919|Aberdeen University
13127|30 March 1937|
10396|26 June 1936|Balliol College, Oxford; Trinity College, Cambridge; Columbia University, New York
13129|20 February 1943|University College, London
13130|19 May 1945|Shenstone Training College; Portsmouth Polytechnic
10406|21 January 1938|Stranmillis Teacher Training College, Belfast 1958
12907|27 November 1945|Newnham College, Cambridge
12905|16 May 1957|
12904|19 September 1940|
12903|10 March 1949|Moray House College of Education; Inverness College
12902|11 September 1931|Trinity College, Cambridge
12901|14 March 1928|Ruskin College, Oxford
12910|16 November 1933|
12909|14 April 1935|London Polytechnic
13551|18 April 1924|London School of Economics
13552|5 September 1938|Birmingham University; London University
13549|8 January 1936|Sydney University, Australia
13626|11 September 1929|Mons Officer Cadet School, Aldershot; Balliol College, Oxford
13632|22 July 1931|Trinity College, Cambridge
13554|1 January 1954|Oxford Polytechnic
13546|13 June 1933|London School of Economics
13547|23 June 1932|Trinity Hall, Cambridge
13286|6 May 1943|London University; Graduate School of Business, Columbia University, New York
13285|27 August 1920|
13287|3 May 1932|Trinity College, Cambridge
13290|20 October 1926|New College, Oxford
13289|6 April 1935|
13276|26 November 1937|London School of Economics
13043|22 September 1924|King's College, Cambridge
13044|16 May 1934|Oriel College, Oxford
13045|28 June 1959|Van Mildert College, Durham University; King's College, London; Institute of Education, London
10446|5 November 1931|University College of Wales, Aberystwyth; Gonville and Caius College, Cambridge; Gray's Inn, Hocker Senior Exhibitioner
13039|23 March 1928|Ruskin College, Oxford 1949-50; St Catherine's College, Oxford; Department of Education, Manchester University
13040|24 November 1922|London School of Economics statistics 1943
13042|13 September 1955|University College, Oxford; Brasenose College, Oxford
13705|10 May 1931|St John's College, Cambridge
13704|25 November 1936|St Catharine's College, Cambridge
13703|8 August 1926|Magdalen College, Oxford; All Souls College, Oxford
13702|14 February 1953|St Catherine's College, Oxford
13709|6 August 1944|Van Mildert College, Durham; Linacre College, Oxford; Ripon Hall, Oxford
13708|29 August 1937|Trinity College, Oxford
13689|25 January 1933|Liverpool University; Trinity Hall, Cambridge
13706|16 October 1941|The Royal Academy of Music
13701|27 November 1929|RMA, Sandhurst
13710|21 March 1923|
13439|23 June 1949|Bristol University
13438|18 February 1926|Magdalen College, Oxford
13435|21 February 1954|Bristol University
13436|3 November 1954|University College, London
13433|25 November 1923|Emmanuel College, Cambridge
13434|21 August 1954|St Anne's College, Oxford; Bryn Mawr College, Pennsylvania University, USA
13441|5 March 1951|Sheffield University; University of Pennsylvania
13442|10 January 1947|University and Nuffield Colleges, Oxford
13165|3 February 1938|University College, Dublin
13167|23 August 1941|Somerville College, Oxford; Harvard University
13166|28 February 1938|Sorbonne
13161|26 July 1930|Royal Academy of Dramatic Art
13163|24 March 1945|Catford College
13162|2 July 1938|Sidney Sussex College, Cambridge; St Thomas's Hospital, London 1956-61
13169|2 November 1934|Oxford University 1957, MA; Princeton University, USA
13168|2 June 1936|RMA, Sandhurst; Selwyn College, Cambridge; Cuddesdon College, Oxford
12945|8 October 1951|Edinburgh University
12946|20 July 1935|Worcester College, Oxford
12947|4 January 1935|Bombay University; London University
12949|1 September 1931|Emmanuel College, Cambridge
12951|11 May 1938|St Andrews University
12937|7 June 1940|MS Baroda University, India
12938|17 July 1945|Sidney Sussex College, Cambridge
13603|18 February 1931|Punjab University; Massachusetts Institute of Technology
13602|20 July 1942|
13601|3 October 1947|Tours University, France; Royal Agricultural College, Cirencester
10475|10 June 1934|Plater Hall, Oxford University
13009|15 October 1931|Girton College, Cambridge 1952, MA
13597|19 March 1931|London School of Economics; Princeton University, USA
13594|15 March 1939|Trinity Hall, Cambridge
12943|21 January 1938|King's College, Cambridge
13425|5 September 1933|Jesus College, Cambridge
13424|4 January 1940|Bristol University
13427|19 March 1945|King's College, London; Hull University
13426|18 April 1923|Girton College, Cambridge
13429|27 March 1925|
12916|27 October 1958|University College, Cardiff; Imperial College, London
13695|6 June 1941|New College, Oxford
13071|29 June 1948|Leeds University; Glasgow University
13693|11 October 1927|Pembroke College, Cambridge
13694|8 December 1923|University College of Wales, Aberystwyth
13699|25 February 1941|City and Guilds 1958-62
13697|25 March 1925|Christ Church, Oxford
13698|12 July 1920|University College, London; Yale University
10495|4 October 1936|Magdalen College, Oxford
13691|12 July 1936|Glasgow University; Graduate Institute for International Affairs, Geneva 1967-68
13038|22 June 1938|
13037|27 January 1939|Le Manoir, Lausanne, Switzerland; Florence University; University College, London; London School of Economics
13244|12 June 1943|Open Scholar Worcester College, Oxford
13033|6 June 1928|Christ's College, Cambridge; University College Hospital, London
13032|19 July 1937|Christ Church, Oxford
13031|18 July 1967|Newcastle University
13291|14 July 1928|Balliol College, Oxford
12967|17 February 1930|
12970|25 July 1937|St John's College, Cambridge; British School of Archaeology, Athens
13277|8 July 1960|Liverpool University
13279|28 May 1932|Magdalen College, Oxford
13280|13 December 1937|Jesus College, Cambridge; University of Paris (Sorbonne)
13281|30 May 1932|Pembroke College, Oxford
13401|24 February 1938|Stockwell College; Wesley Deaconess College; Wesley House, Cambridge
13332|27 January 1924|
13331|10 July 1930|University College, Oxford
10504|12 April 1946|Dundee University
13328|18 September 1944|Glasgow University; New College, Oxford
13327|28 October 1928|Magdalen College, Oxford
13330|30 June 1942|Belfast Institute of Technology; The Open University
13329|23 July 1933|Architectural Association; Yale University; RIBA
10511|5 June 1941|Handsworth Technical College 1957-60; Aston University; Warwick University
13005|10 September 1935|Magdalen College, Oxford; University of Chicago
13006|31 March 1958|Bristol University; Cambridge University
13592|12 March 1954|RMA, Sandhurst; Royal Agricultural College, Cirencester
13588|4 February 1949|Magdalene College, Cambridge
13589|21 June 1946|London School of Economics
13022|2 November 1927|Worcester College, Oxford
13026|24 October 1940|King's College, Cambridge; Columbia University, New York
13625|16 May 1957|
13624|18 May 1929|Fitzwilliam College, Cambridge; Christ Church, Oxford; Yale University, USA
13628|1 October 1942|Trinity College, Oxford; Cuddesdon Theological College
12942|18 October 1930|
12941|31 May 1927|
12912|30 April 1933|Bradford Technical College; Scottish College of Textiles
13633|11 April 1943|Trinity College, Cambridge; OU certificate in European studies 1973
13145|20 March 1936|Brasenose College, Oxford
13146|12 May 1943|
13141|19 August 1955|London University
13142|2 October 1934|Cape Town University; Trinity College, Cambridge
13143|10 August 1957|University of East Anglia
13144|3 May 1930|
13181|24 March 1940|Christ Church, Oxford
13182|31 July 1942|Balliol College, Oxford; Edinburgh University
13184|27 October 1937|
13183|15 January 1946|Durham University; University College of Wales, Swansea; Aberdeen University
13186|19 February 1943|
13185|21 November 1938|Newnham College, Cambridge
13188|11 February 1923|Florence
13187|9 October 1920|
10535|13 September 1923|London University
13191|25 December 1932|London School of Economics
13152|18 Dec 1952|
13455|16 March 1942|
13456|20 July 1940|School of Navigation, Southampton University; Sydney Technical College
13462||
13459||
13460|2 April 1945|Somerset Farm Institute; Hadlow College of Agriculture and Horticulture
13463|25 April 1939|Jesus College, Oxford
13464|20 July 1927|
13654|14 June 1937|London School of Economics
13324|4 June 1940|Glasgow University
13326|24 July 1945|London School of Economics; Garnett College, London University; Salford University
13657|7 March 1930|Jesus College, Cambridge
13658|23 June 1926|Edinburgh University; Cambridge University
13337|31 March 1938|Edinburgh University
13338|27 December 1934|Guildhall School of Music
13385|25 September 1941|Bristol University
13384|26 May 1936|Sidney Sussex College, Cambridge
13387|19 July 1945|King's College, Cambridge
13386|10 August 1935|Jesus College, Cambridge
13389|15 August 1932|University of Stellenbosch, South Africa; University College, Oxford
13557|4 May 1926|
13630|7 September 1942|
13629|1 November 1914|Chelsea School of Art
13203|22 February 1960|University of East Anglia 1978-82; University of Aix-en-Provence 1981
13204|25 February 1941|Aberdeen University; Corpus Christi College, Cambridge
13205|14 December 1938|RMA, Sandhurst
13206|14 April 1951|Girton College, Cambridge
13207|30 March 1934|Trinity College, Cambridge
13208|18 October 1928|Balliol College, Oxford
13209|10 June 1929|
13194|21 September 1952|Keele University; Gray's Inn, Inns of Court School of Law
13195|29 March 1931|
12978|3 March 1920|St John's College, Cambridge
10592|12 February 1938|St. Catharine's College, Cambridge
12976|7 November 1927|St Catharine's College, Cambridge
12975|13 October 1925|Somerville College, Oxford
12974|13 March 1937|Peterhouse, Cambridge
12972|19 October 1937|School of Management, Bath University; INSEAD (AMP) 1987
12971|21 October 1931|Queens' College, Cambridge; Sorbonne, Paris
12935|20 December 1935|Lady Margaret Hall, Oxford University
13543|16 October 1952|London School of Economics
13544|17 May 1924|Birmingham College of Technology; London University
13541|1 August 1939|Co-operative College, Loughborough; Brunel University; Warwick University
13542|30 November 1943|
13539|11 October 1928|Manchester University
13540|31 March 1941|Princeton University, USA
13538|23 October 1922|
13536|23 February 1937|Gonville and Caius College, Cambridge
13272|22 March 1934|Manchester University
13271|18 September 1927|
13274|17 July 1959|Polytechnic of North London
13273|9 January 1942|Trinity College, Cambridge
13267|23 August 1931|Royal Military College of Science
13270|27 January 1931|
13264|2 August 1929|Hertford College, Oxford
13263|24 December 1932|Queen's University, Belfast
13114|22 June 1932|
13115|15 August 1946|Corpus Christi College, Oxford; Harvard University 1969-70
13117|17 March 1938|Trinity College, Cambridge
13110|25 March 1932|
13112|12 March 1941|King's College, Cambridge; Cornell University, USA; Nuffield College, Oxford
13113|12 April 1943|Liverpool University; Manchester Polytechnic
13119|8 December 1938|King's College, Cambridge
13120|16 September 1922|Medical School, King's College, Newcastle upon Tyne (Durham University)
12896|8 September 1940|University of California, Berkeley
12895|14 April 1924|Lady Margaret Hall, Oxford
12894|16 July 1945|Bedford College, London University
12893|1 May 1949|Heriot-Watt University, Edinburgh
12900|3 February 1941|Jesus College, Cambridge
12899|31 October 1949|
12897|13 April 1927|Queens' College, Cambridge
12888|13 September 1919|Vienna University
12957|20 Feb 1936|Girton College, Cambridge; Bryn Mawr College, USA; Harvard University, USA
12958|15 June 1943|St John's College, Cambridge
12961|31 October 1940|Plymouth University
12962|6 May 1946|Manchester University
12959|27 July 1930|Somerville College, Oxford; Columbia University, New York
12960|9 February 1933|Christ Church, Oxford; London School of Economics
13617|8 May 1934|Exeter College, Oxford
13072|14 September 1938|New College, Oxford
13616|11 October 1942|
13619|14 February 1935|Keble College, Oxford; London University
13618|15 March 1943|King's College, Cambridge; Cuddesdon Theological College
13621|28 January 1932|Trinity College, Oxford; Brasenose College, Oxford
13620|15 July 1940|London Hospital Medical College, London University
13623|11 November 1927|
13622|9 November 1935|Trinity College, Cambridge; Stanford University, California, USA
13615|2 May 1933|University College, London
13614|25 April 1940|Leeds University
13025|28 June 1931|Merton College, Oxford
13023|27 February 1932|University College, London
13030|8 April 1948|Edinburgh University; Strathclyde University; DipHSM 1974
13294|5 March 1960|Aston University Production engineering 1982, PhD robotics 1985
13197|21 November 1931|
13196|6 June 1940|IIT, Kharagpur; Birmingham University
13548|9 March 1955|London School of Economics; University of Kent
13545|10 November 1943|Bedford College, London; Lancaster University
13201|22 April 1941|
13200|29 Jun 1940|
13199|9 February 1946|Durham University
13198||
12845|20 March 1959|Exeter College, Oxford
13558|14 Nov 1941|
13481|5 October 1944|University of London economics 1970
13482|16 January 1947|Manchester University; University College, London
13483|18 January 1938|Hull University; London School of Economics; University of Cambridge
10554|12 February 1942|
13477|23 October 1935|University College of North Wales; Handsworth Methodist College
13478|20 September 1938|Punjab University
13479|20 October 1947|
13480|30 August 1961|Bedford College, London
13475|22 August 1937|North East London Polytechnic
10425|5 May 1936|University College, Oxford
13055|27 February 1950|Newnham College, Cambridge; Leo Baeck College, London
13056|5 January 1944|
13057|24 July 1946|Bristol University
13058|26 Jun 1961|
13051|17 May 1939|Pembroke College, Cambridge
13052|26 April 1948|St Andrews University; Barking Regional College of Technology
13053|30 March 1950|East London College; Sussex University; London School of Economics; London Business School
13054|17 September 1938|Melbourne University, Australia; Gonville and Caius College, Cambridge
13048|1 June 1951|New College of Speech and Drama; Middlesex Polytechnic/University
10516|23 January 1940|King's College, London
12838|20 October 1957|University College, London
12837|15 February 1942|University College of Wales, Cardiff; Fitzwilliam College, Cambridge; School of Oriental and African Studies, London University
12836|17 January 1943|University College, London; College of Air Training, Hamble
12835|22 December 1942|Leeds University; Columbia University, New York, USA
12842|28 June 1934|Pembroke College, Oxford; Chicago University Law School
12841|9 April 1937|Worcester College, Oxford
12840|31 January 1945|Girton College, Cambridge
12839|30 October 1943|Essex University; King's College, Cambridge
12844|19 January 1951|Lancaster University; Oxford University; Cuddesdon Theological College, Oxford
12843|20 May 1943|Brasenose College, Oxford; London Business School
13450|14 April 1942|
13447|24 November 1949|Oxford University
13445|15 June 1932|
13443|22 February 1942|Pembroke College, Oxford
13444|18 April 1944|University College, London; Lady Margaret Hall, Oxford
13452|20 August 1955|London University
13453|31 December 1946|Selwyn College, Cambridge; Ripon Hall, Oxford
13177|12 Mar 1951|Trinity College, Cambridge
13176|12 May 1944|Balliol College, Oxford Oxford
13171|28 March 1942|University College of Wales, Cardiff
13170|30 Jul 1939|
13173|30 June 1957|
13172|20 Apr 1931|Magdalen College, Oxford
13179|14 Apr 1940|Nottingham University; St Stephen's House; Linacre College, Oxford
13178|22 February 1963|Keble College, Oxford; Christ Church, Oxford
13149|6 November 1934|Corpus Christi College, Cambridge
13150|21 Oct 1942|Leicester University; Southampton University
13151|2 December 1956|Lincoln College, Oxford
10345|22 April 1946|Heriot-Watt University
10584|2 July 1947|Bradford University; Sheffield University
10464|6 January 1945|Heriot-Watt University; Moray House College of Education, Edinburgh
10612|29 October 1941|Exeter College, Oxford
10445|17 June 1952|Coventry College of Education
10291|11 June 1944|King's College, Cambridge
10207|25 June 1937|Oxford University
10101|9 July 1942|Portsmouth Polytechnic; Portsmouth Naval College; Graduate, Institute of Mechanical Engineers
10599|19 February 1941|University College, London
10211|21 January 1942|Edinburgh University
10255|30 December 1941|
12928|18 August 1928|Trinity College, Cambridge
10325|30 March 1948|
10536|22 January 1940|St Hilda's College, Oxford
10374|27 Mar 1939|Christ Church, Oxford; College of Law
12933||Birmingham University; Filtzwilliam College, Cambridge; Ridley Hall, Cambridge
10607||
13583|25 February 1947|St Andrews University; Edinburgh University
10058|12 March 1948|Essex University; London School of Economics
10424|26 July 1940|Queen's University, Belfast; Michigan University, USA; London University
10110|26 February 1949|Queens College, St Andrews University; Edinburgh University
10556|7 May 1939|Newbattle Abbey Adult Education College; Strathclyde University; Southampton University
10547|24 July 1951|Pembroke College, Cambridge; Harvard University
10003|27 December 1947|
13577|29 April 1942|
10011|17 June 1939|University College of Wales, Swansea; Inns of Court School of Law 1966-69
10135|5 May 1942|London School of Economics; Inns of Court School of Law 1989-90; Open University
10234|4 Jul 1943|King's College, Cambridge
13683||
10146|4 August 1939|Bede College, Durham University
13321|6 June 1943|University College, Oxford
13320|5 October 1955|Gonville and Caius College, Cambridge
13323|23 June 1942|Trinity College, Cambridge
13322|29 April 1943|St Anne's College, Oxford; Brandess University, USA
13315|8 December 1958|St Hugh's College, Oxford
13714|10 June 1949|Makere Iniversity, Uganda; Diploma in legal practice, Uganda 1972; Selwyn College, Cambridge; Ridley Hall, Cambridge
13716|21 January 1945|Christ's College, Cambridge
13718||
13717||
10136||
13720||
13721||
13724||
13723||
13725||
13727||
13728||
13726||
13730||
13729||
13731||
13732||
13734||
13733||
13737||
13740||
13739||
13876||
13877||
10059||
13880||
13882||
13878||Queen's University, Belfast
13881||
13879||
13883||
13884||
13885||
13886||
13738||
13890||
13920||
13919||
13922||
13921||
13923||
13924||
13925||
13926||
13929||
13928||
13931||
13932||
13937||
13936||
13939||
13938||
13940||
10605||
14126||
14125||
14127||
14129||
14130||
14132||
14133||
14134||
14135||
13261||
14136||
14138||
10412||
14139||
14140||
14143||
14144||
14145||
14147||
24686||
24685||
24687||
24688||
24689||
13930||
24690||
24693||
24692||
10420||
24694||
24695||
24696||
24700||
24699||
24698||
24706||
24705||
24704||
